module custom_or(input a,b,output w);
    c1 c(1'b0 , 1'b0 , 1'b0 , 1'b1 , 1'b1 ,1'b0 , a , b, w) ;
endmodule