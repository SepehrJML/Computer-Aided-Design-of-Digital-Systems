module custom_and(input a,b,output w);
    c1 c(1'b0 , b , a , 1'b0 , 1'b0 ,1'b0 , 1'b0 , 1'b0, w) ;
endmodule