module custom_not(input a,output w);
    c1 c( 1'b1 , 1'b0 , a , 1'b0 , 1'b0 ,1'b0 , 1'b0 , 1'b0, w) ;
endmodule